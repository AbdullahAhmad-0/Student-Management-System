Demo:210.297.mm
a:210.297.mm